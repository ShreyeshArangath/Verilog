module greater_than(A,B,F);

input[1:0] //Since we want a two bit number. If we needed an 8 bit number: input[7:0]

endmodule